/*
Copyright by Henry Ko and Nicola Nicolici
Developed for the Digital Systems Design course (COE3DQ4)
Department of Electrical and Computer Engineering
McMaster University
Ontario, Canada
*/

`timescale 1ns/100ps
`default_nettype none

module SRAM_BIST (
	input logic Clock,
	input logic Resetn,
	input logic BIST_start,
	
	output logic [17:0] BIST_address,
	output logic [15:0] BIST_write_data,
	output logic BIST_we_n,
	input logic [15:0] BIST_read_data,
	
	output logic BIST_finish,
	output logic BIST_mismatch
);

enum logic [2:0] {
	S_IDLE,
	S_DELAY_1,
	S_DELAY_2,
	S_WRITE_CYCLE,
	S_READ_CYCLE,
	S_DELAY_3,
	S_DELAY_4
} BIST_state;

logic BIST_start_buf;

// no need to keep the data that is written into the memory (or comapared against while reading) in a separate register
assign BIST_write_data = BIST_address[15:0];

// mode is 0 for the first burst and mode is 1 for the second burst
logic BIST_mode;

// The BIST engine
always_ff @ (posedge Clock or negedge Resetn) begin
	if (Resetn == 1'b0) begin
		BIST_state <= S_IDLE;
		BIST_mismatch <= 1'b0;
		BIST_finish <= 1'b0;
		BIST_address <= 18'd0;
		BIST_we_n <= 1'b1;		
		BIST_start_buf <= 1'b0;
		BIST_mode <= 1'b0;
	end else begin
		BIST_start_buf <= BIST_start;		
		case (BIST_state)
		S_IDLE: begin
			if (BIST_start & ~BIST_start_buf) begin
				// Start the BIST engine
				BIST_address <= 18'h1FFFF; // jump at the end of the first segment
				BIST_we_n <= 1'b0;
				BIST_mismatch <= 1'b0;
				BIST_finish <= 1'b0;
				BIST_mode <= 1'b0;
				BIST_state <= S_WRITE_CYCLE;
			end else begin
				BIST_address <= 18'd0;
				BIST_we_n <= 1'b1;
				BIST_finish <= 1'b1;
			end
		end
		S_DELAY_1: begin
			BIST_address <= (BIST_mode == 1'b0) ? BIST_address + 18'd1 : BIST_address - 18'd1;
			BIST_state <= S_DELAY_2;
		end
		S_DELAY_2: begin
			BIST_address <= (BIST_mode == 1'b0) ? BIST_address + 18'd1 : BIST_address - 18'd1;
			BIST_state <= S_READ_CYCLE;
		end
		S_WRITE_CYCLE: begin
			if (BIST_mode == 1'b0) begin
				if (BIST_address == 18'd0) begin
					BIST_we_n <= 1'b1;
 					BIST_state <= S_DELAY_1;
 				end
				else
					BIST_address <= BIST_address - 18'd1;
			end else begin
				if (BIST_address == 18'h3FFFF) begin
					BIST_we_n <= 1'b1;
 					BIST_state <= S_DELAY_1;
 				end
				else
					BIST_address <= BIST_address + 18'd1;
			end
		end
		S_READ_CYCLE: begin
			if (BIST_mode == 1'b0) begin
				if (BIST_read_data != (BIST_write_data - 16'd2)) 
					BIST_mismatch <= 1'b1;
				BIST_address <= BIST_address + 18'd1;								
				if (BIST_address == 18'h1FFFF) begin
					BIST_we_n <= 1'b0;
					BIST_state <= S_DELAY_3;
				end
			end else begin
				if (BIST_read_data != (BIST_write_data + 16'd2)) 
					BIST_mismatch <= 1'b1;
				BIST_address <= BIST_address - 18'd1;								
				if (BIST_address == 18'h20000) begin
					BIST_state <= S_DELAY_3;
				end
			end
		end
		S_DELAY_3: begin
			if (BIST_read_data != (BIST_write_data + ((BIST_mode == 1'b0) ? -16'd2 : 16'd2))) 
				BIST_mismatch <= 1'b1;
			BIST_address <= (BIST_mode == 1'b0) ? BIST_address + 18'd1 : BIST_address - 18'd1;
			BIST_state <= S_DELAY_4;
		end
		S_DELAY_4: begin
			if (BIST_read_data != (BIST_write_data + ((BIST_mode == 1'b0) ? -16'd2 : 16'd2))) 
				BIST_mismatch <= 1'b1;
			BIST_address <= (BIST_mode == 1'b0) ? BIST_address + 18'd1 : 18'd0;
			if (BIST_mode == 1'b0) begin
				BIST_mode <= 1'b1;
				BIST_state <= S_WRITE_CYCLE;
			end else begin
				BIST_mode <= 1'b0;
				BIST_finish <= 1'b1;
				BIST_state <= S_IDLE;
			end
		end
		default: BIST_state <= S_IDLE;
		endcase
	end
end

endmodule
